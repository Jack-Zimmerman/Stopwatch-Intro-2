module tb_timer();
	localparam FREQUENCY = 10_000_000;
	localparam MAX_SECONDS = 10;

endmodule
